module top_module(
    input a,
    input b,
    input c,
    output wire out  ); 
    or or1(out,a,b,c);
endmodule
