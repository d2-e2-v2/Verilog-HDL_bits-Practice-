module top_module(
    input [31:0] a,
    input [31:0] b,
    output [31:0] sum
);
    wire cin,cout;
    add16 k1(.a(a[15:0]),.b(b[15:0]),.sum(sum[15:0]),.cin(0),.cout(cin));
    add16 k2(.a(a[31:16]),.b(b[31:16]),.cin(cin),.cout(cout),.sum(sum[31:16]));

endmodule
