module top_module ( input x, input y, output z );
    xnor nor1(z,x,y);
endmodule
